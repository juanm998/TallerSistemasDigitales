package my_pkg is
    type t_estado is (E_R1_V2, E_R1_A2, E_A1_R2, E_V1_R2, E_R2_A1, E_A2_R1);
end my_pkg;